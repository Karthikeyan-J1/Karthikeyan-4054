1.STEP ONE:
module top_module( output one );

// Insert your code here
    assign one = 1;

endmodule

2.ZERO:
module top_module(
    output zero
);// Module body starts after semicolon
assign zero=0;
endmodule
